/* TinyQV: A RISC-V core designed to use minimal area.
  
   This memory controller plumbs the outputs from the CPU into the Flash and RAM controllers
 */

module tinyqv_mem_ctrl (
    input clk,
    input rstn,

    input [23:1] instr_addr,
    input        instr_jump,
    input        instr_fetch_stall,

    output       instr_ready,

    input [24:0] data_addr,
    input [1:0]  data_write_n, // 11 = no write, 00 = 8-bits, 01 = 16-bits, 10 = 32-bits
    input [1:0]  data_read_n,  // 11 = no read,  00 = 8-bits, 01 = 16-bits, 10 = 32-bits
    input [31:0] data_to_write,

    input        data_continue, // Whether another read/write at the next address will immediately follow this one

    output         data_ready,  // Transaction complete/data request can be modified.
    output  [31:0] data_from_read,

    // External SPI interface
    input      [3:0] spi_data_in,
    output     [3:0] spi_data_out,
    output     [3:0] spi_data_oe,
    output           spi_clk_out,
    output           spi_flash_select,
    output           spi_ram_a_select,
    output           spi_ram_b_select,

    output        debug_stall_txn,
    output        debug_stop_txn
);

    // Combinational
    reg start_instr;
    reg start_read;
    reg start_write;
    reg stop_txn;
    reg continue_txn;
    reg [1:0] data_txn_n;
    reg [1:0] data_txn_len;

    reg qspi_write_done;
    wire qspi_busy;
    reg instr_active;
    reg instr_fetch_restart;

    wire is_instr = instr_active || start_instr;
    wire [1:0] txn_len = is_instr ? 2'b11 : data_txn_len;
    wire [24:0] addr_in = is_instr ? {1'b0, instr_addr, 1'b0} : data_addr[24:0];
    reg [31:0] qspi_data_buf;
    reg [1:0] qspi_data_byte_idx;
    wire qspi_data_req;
    wire qspi_data_ready;
    wire [7:0] qspi_data_out;

    // Only stall on the last byte of an instruction
    wire stall_txn = instr_active && instr_fetch_stall && !instr_ready && qspi_data_byte_idx == 2'b11;
    reg data_stall;

    always @(*) begin
        start_instr = 0;
        start_read = 0;
        start_write = 0;
        stop_txn = 0;
        data_txn_n = data_write_n & data_read_n;

        if (qspi_busy || qspi_write_done) begin
            // A transaction is running
            if (instr_active) begin
                if (instr_fetch_restart || data_txn_n != 2'b11) begin
                    // Stop immediately on restart or data txn
                    stop_txn = 1;
                end
            end else if ((qspi_data_ready || qspi_data_req) && qspi_data_byte_idx == data_txn_len && !continue_txn) begin
                // Data transaction is complete
                stop_txn = 1;
            end
        end else begin
            // No transaction, start one
            if (data_read_n != 2'b11)
                start_read = 1;
            else if (data_write_n != 2'b11)
                start_write = 1;
            else if (instr_fetch_restart)
                start_instr = 1;
        end
    end

    // State
    always @(posedge clk) begin
        if (!rstn || stop_txn) begin
            instr_active <= 0;
        end else begin
            instr_active <= qspi_busy ? instr_active : start_instr;
        end
    end

    wire [1:0] write_qspi_data_byte_idx = qspi_data_byte_idx + (qspi_data_req ? 2'b01 : 2'b00);
    qspi_controller q_ctrl(
        .clk(clk),
        .rstn(rstn),

        .spi_data_in(spi_data_in),
        .spi_data_out(spi_data_out),
        .spi_data_oe(spi_data_oe),
        .spi_clk_out(spi_clk_out),

        .spi_flash_select(spi_flash_select),
        .spi_ram_a_select(spi_ram_a_select),
        .spi_ram_b_select(spi_ram_b_select),

        .addr_in(addr_in),
        .data_in(qspi_data_buf[{write_qspi_data_byte_idx,3'b000} +:8]),
        .start_read(start_read || start_instr),
        .start_write(start_write),
        .stall_txn(stall_txn || data_stall),
        .stop_txn(stop_txn),

        .data_out(qspi_data_out),
        .data_req(qspi_data_req),
        .data_ready(qspi_data_ready),
        .busy(qspi_busy)
    );

    always @(posedge clk) begin
        if (!rstn) begin
            instr_fetch_restart <= 1'b0;
        end else begin
            instr_fetch_restart <= start_instr ? 1'b0 : stop_txn | !instr_active | instr_jump;
        end
    end

    always @(posedge clk) begin
        if (!rstn || start_instr || start_read || start_write) begin
            qspi_data_byte_idx <= 2'b00;
        end else begin
            if (qspi_data_ready || qspi_data_req) begin
                qspi_data_byte_idx <= qspi_data_byte_idx + 2'b01;

                if (qspi_data_byte_idx == txn_len) begin
                    qspi_data_byte_idx <= 0;
                end
            end
        end
    end

    always @(posedge clk) begin
        if (qspi_data_ready) begin
            qspi_data_buf[{qspi_data_byte_idx,3'b000} +:8] <= qspi_data_out;
        end else if (data_write_n != 2'b11 && (data_stall || start_write)) begin
            qspi_data_buf <= data_to_write;
        end
    end

    assign instr_ready = instr_active && qspi_data_ready && qspi_data_byte_idx == 2'b11;

    always @(posedge clk) begin
        qspi_write_done <= qspi_data_req && qspi_data_byte_idx == data_txn_len;
    end

    always @(posedge clk) begin
        if (!rstn)
            data_txn_len <= 2'b11;
        else if (start_read || start_write) begin
            data_txn_len <= {data_txn_n[1], data_txn_n[1] | data_txn_n[0]};  // 0, 1 or 3 for 1, 2 or 4 byte txn
        end
    end

    always @(posedge clk) begin
        if (!rstn) begin
            continue_txn <= 0;
        end else begin
            if (continue_txn) begin
                if ((qspi_data_req && qspi_data_byte_idx + 2'b01 == data_txn_len) ||
                    (qspi_data_ready && qspi_data_byte_idx == data_txn_len))
                begin
                    data_stall <= 1;
                end else if (data_stall && qspi_data_byte_idx == 2'b00 && ((data_read_n != 2'b11 && !data_ready) || data_write_n != 2'b11)) begin
                    data_stall <= 0;
                    continue_txn <= data_continue;
                end
            end else begin
                data_stall <= 0;
                if (start_write || start_read) begin
                    continue_txn <= data_continue;
                end
            end
        end
    end

    assign data_ready = !instr_active && ((qspi_data_ready && qspi_data_byte_idx == data_txn_len) || (data_write_n != 2'b11 && ((data_stall && qspi_data_byte_idx == 2'b00) || (data_continue ? start_write : qspi_write_done))));
    assign data_from_read = (qspi_data_ready && qspi_data_byte_idx == txn_len) ? 
      ({qspi_data_out, qspi_data_buf[23:16],
        txn_len == 2'b01 ? qspi_data_out : qspi_data_buf[15:8],
        txn_len == 2'b00 ? qspi_data_out : qspi_data_buf[7:0]}) : qspi_data_buf;

    assign debug_stall_txn = stall_txn;
    assign debug_stop_txn = stop_txn;

endmodule
